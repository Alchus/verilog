/*
HelloWorld.v
By Thomas Sowders
CONTENTS:
module helloworld - Displays a cheerful message.
*/

/*
MODULE helloworld
By Thomas Sowders
Description:
	Prints a cheerful message.
Arguments:
	(none)
*/
module helloworld;
	initial
	//Display the text "Hello World"
	$display("Hello World \n Thomas Sowders");
endmodule