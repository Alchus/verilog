module Test ();
initial
 $display("Hello world");

endmodule